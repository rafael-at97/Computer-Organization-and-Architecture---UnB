cte10_inst : cte10 PORT MAP (
		result	 => result_sig
	);
