cte22_inst : cte22 PORT MAP (
		result	 => result_sig
	);
