shiftl2_inst : shiftl2 PORT MAP (
		data	 => data_sig,
		distance	 => distance_sig,
		result	 => result_sig
	);
