ULAaddcte_inst : ULAaddcte PORT MAP (
		result	 => result_sig
	);
