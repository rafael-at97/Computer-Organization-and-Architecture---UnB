ula_multu_inst : ula_multu PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		result	 => result_sig
	);
