shiftarithmetic_inst : shiftarithmetic PORT MAP (
		data	 => data_sig,
		distance	 => distance_sig,
		result	 => result_sig
	);
