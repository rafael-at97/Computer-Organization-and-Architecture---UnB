ADD4_inst : ADD4 PORT MAP (
		dataa	 => dataa_sig,
		result	 => result_sig
	);
